`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/06/2020 02:50:06 PM
// Design Name: 
// Module Name: rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module rom
(
   input i_clk,
   input i_ce,
   input i_rst,
   output signed [15:0] o_data
);

(*rom_style = "block" *) reg signed [15:0] s;
reg [9:0] addr;

assign o_data = s;

always @(posedge i_clk) begin
    if (i_rst)
        addr <= 0;
    else if (i_ce)
        addr <= addr + 1'b1;
end

always @(posedge i_clk) begin
    if (i_ce)
        case (addr)
            10'd0: s <= 16'd9830;
            10'd1: s <= 16'd24018;
            10'd2: s <= -16'd20394;
            10'd3: s <= 16'd12457;
            10'd4: s <= -16'd8514;
            10'd5: s <= -16'd25966;
            10'd6: s <= 16'd15986;
            10'd7: s <= -16'd17503;
            10'd8: s <= 16'd4915;
            10'd9: s <= 16'd25301;
            10'd10: s <= -16'd13443;
            10'd11: s <= 16'd22203;
            10'd12: s <= -16'd1;
            10'd13: s <= -16'd22204;
            10'd14: s <= 16'd13442;
            10'd15: s <= -16'd25302;
            10'd16: s <= -16'd4916;
            10'd17: s <= 16'd17502;
            10'd18: s <= -16'd15987;
            10'd19: s <= 16'd25965;
            10'd20: s <= 16'd8513;
            10'd21: s <= -16'd12458;
            10'd22: s <= 16'd20393;
            10'd23: s <= -16'd24019;
            10'd24: s <= -16'd9831;
            10'd25: s <= 16'd8420;
            10'd26: s <= -16'd25482;
            10'd27: s <= 16'd19981;
            10'd28: s <= 16'd8513;
            10'd29: s <= -16'd6474;
            10'd30: s <= 16'd29888;
            10'd31: s <= -16'd14937;
            10'd32: s <= -16'd4916;
            10'd33: s <= 16'd7137;
            10'd34: s <= -16'd32434;
            10'd35: s <= 16'd10234;
            10'd36: s <= -16'd1;
            10'd37: s <= -16'd10235;
            10'd38: s <= 16'd32433;
            10'd39: s <= -16'd7138;
            10'd40: s <= 16'd4915;
            10'd41: s <= 16'd14936;
            10'd42: s <= -16'd29889;
            10'd43: s <= 16'd6473;
            10'd44: s <= -16'd8514;
            10'd45: s <= -16'd19982;
            10'd46: s <= 16'd25481;
            10'd47: s <= -16'd8421;
            10'd48: s <= 16'd9830;
            10'd49: s <= 16'd24018;
            10'd50: s <= -16'd20394;
            10'd51: s <= 16'd12457;
            10'd52: s <= -16'd8514;
            10'd53: s <= -16'd25966;
            10'd54: s <= 16'd15986;
            10'd55: s <= -16'd17503;
            10'd56: s <= 16'd4915;
            10'd57: s <= 16'd25301;
            10'd58: s <= -16'd13443;
            10'd59: s <= 16'd22203;
            10'd60: s <= 16'd0;
            10'd61: s <= -16'd22204;
            10'd62: s <= 16'd13442;
            10'd63: s <= -16'd25302;
            10'd64: s <= -16'd4916;
            10'd65: s <= 16'd17502;
            10'd66: s <= -16'd15987;
            10'd67: s <= 16'd25965;
            10'd68: s <= 16'd8513;
            10'd69: s <= -16'd12458;
            10'd70: s <= 16'd20393;
            10'd71: s <= -16'd24019;
            10'd72: s <= -16'd9831;
            10'd73: s <= 16'd8420;
            10'd74: s <= -16'd25482;
            10'd75: s <= 16'd19981;
            10'd76: s <= 16'd8513;
            10'd77: s <= -16'd6474;
            10'd78: s <= 16'd29888;
            10'd79: s <= -16'd14937;
            10'd80: s <= -16'd4916;
            10'd81: s <= 16'd7137;
            10'd82: s <= -16'd32434;
            10'd83: s <= 16'd10234;
            10'd84: s <= -16'd1;
            10'd85: s <= -16'd10235;
            10'd86: s <= 16'd32433;
            10'd87: s <= -16'd7138;
            10'd88: s <= 16'd4915;
            10'd89: s <= 16'd14936;
            10'd90: s <= -16'd29889;
            10'd91: s <= 16'd6473;
            10'd92: s <= -16'd8514;
            10'd93: s <= -16'd19982;
            10'd94: s <= 16'd25481;
            10'd95: s <= -16'd8421;
            10'd96: s <= 16'd9830;
            10'd97: s <= 16'd24018;
            10'd98: s <= -16'd20394;
            10'd99: s <= 16'd12457;
            10'd100: s <= -16'd8514;
            10'd101: s <= -16'd25966;
            10'd102: s <= 16'd15986;
            10'd103: s <= -16'd17503;
            10'd104: s <= 16'd4915;
            10'd105: s <= 16'd25301;
            10'd106: s <= -16'd13443;
            10'd107: s <= 16'd22203;
            10'd108: s <= 16'd0;
            10'd109: s <= -16'd22204;
            10'd110: s <= 16'd13442;
            10'd111: s <= -16'd25302;
            10'd112: s <= -16'd4916;
            10'd113: s <= 16'd17502;
            10'd114: s <= -16'd15987;
            10'd115: s <= 16'd25965;
            10'd116: s <= 16'd8513;
            10'd117: s <= -16'd12458;
            10'd118: s <= 16'd20393;
            10'd119: s <= -16'd24019;
            10'd120: s <= -16'd9831;
            10'd121: s <= 16'd8420;
            10'd122: s <= -16'd25482;
            10'd123: s <= 16'd19981;
            10'd124: s <= 16'd8513;
            10'd125: s <= -16'd6474;
            10'd126: s <= 16'd29888;
            10'd127: s <= -16'd14937;
            10'd128: s <= -16'd4916;
            10'd129: s <= 16'd7137;
            10'd130: s <= -16'd32434;
            10'd131: s <= 16'd10234;
            10'd132: s <= -16'd1;
            10'd133: s <= -16'd10235;
            10'd134: s <= 16'd32433;
            10'd135: s <= -16'd7138;
            10'd136: s <= 16'd4915;
            10'd137: s <= 16'd14936;
            10'd138: s <= -16'd29889;
            10'd139: s <= 16'd6473;
            10'd140: s <= -16'd8514;
            10'd141: s <= -16'd19982;
            10'd142: s <= 16'd25481;
            10'd143: s <= -16'd8421;
            10'd144: s <= 16'd9830;
            10'd145: s <= 16'd24018;
            10'd146: s <= -16'd20394;
            10'd147: s <= 16'd12457;
            10'd148: s <= -16'd8514;
            10'd149: s <= -16'd25966;
            10'd150: s <= 16'd15986;
            10'd151: s <= -16'd17503;
            10'd152: s <= 16'd4915;
            10'd153: s <= 16'd25301;
            10'd154: s <= -16'd13443;
            10'd155: s <= 16'd22203;
            10'd156: s <= 16'd0;
            10'd157: s <= -16'd22204;
            10'd158: s <= 16'd13442;
            10'd159: s <= -16'd25302;
            10'd160: s <= -16'd4916;
            10'd161: s <= 16'd17502;
            10'd162: s <= -16'd15987;
            10'd163: s <= 16'd25965;
            10'd164: s <= 16'd8513;
            10'd165: s <= -16'd12458;
            10'd166: s <= 16'd20393;
            10'd167: s <= -16'd24019;
            10'd168: s <= -16'd9831;
            10'd169: s <= 16'd8420;
            10'd170: s <= -16'd25482;
            10'd171: s <= 16'd19981;
            10'd172: s <= 16'd8513;
            10'd173: s <= -16'd6474;
            10'd174: s <= 16'd29888;
            10'd175: s <= -16'd14937;
            10'd176: s <= -16'd4916;
            10'd177: s <= 16'd7137;
            10'd178: s <= -16'd32434;
            10'd179: s <= 16'd10234;
            10'd180: s <= 16'd0;
            10'd181: s <= -16'd10235;
            10'd182: s <= 16'd32433;
            10'd183: s <= -16'd7138;
            10'd184: s <= 16'd4915;
            10'd185: s <= 16'd14936;
            10'd186: s <= -16'd29889;
            10'd187: s <= 16'd6473;
            10'd188: s <= -16'd8514;
            10'd189: s <= -16'd19982;
            10'd190: s <= 16'd25481;
            10'd191: s <= -16'd8421;
            10'd192: s <= 16'd9830;
            10'd193: s <= 16'd24018;
            10'd194: s <= -16'd20394;
            10'd195: s <= 16'd12457;
            10'd196: s <= -16'd8514;
            10'd197: s <= -16'd25966;
            10'd198: s <= 16'd15986;
            10'd199: s <= -16'd17503;
            10'd200: s <= 16'd4915;
            10'd201: s <= 16'd25301;
            10'd202: s <= -16'd13443;
            10'd203: s <= 16'd22203;
            10'd204: s <= 16'd0;
            10'd205: s <= -16'd22204;
            10'd206: s <= 16'd13442;
            10'd207: s <= -16'd25302;
            10'd208: s <= -16'd4916;
            10'd209: s <= 16'd17502;
            10'd210: s <= -16'd15987;
            10'd211: s <= 16'd25965;
            10'd212: s <= 16'd8513;
            10'd213: s <= -16'd12458;
            10'd214: s <= 16'd20393;
            10'd215: s <= -16'd24019;
            10'd216: s <= -16'd9831;
            10'd217: s <= 16'd8420;
            10'd218: s <= -16'd25482;
            10'd219: s <= 16'd19981;
            10'd220: s <= 16'd8513;
            10'd221: s <= -16'd6474;
            10'd222: s <= 16'd29888;
            10'd223: s <= -16'd14937;
            10'd224: s <= -16'd4916;
            10'd225: s <= 16'd7137;
            10'd226: s <= -16'd32434;
            10'd227: s <= 16'd10234;
            10'd228: s <= 16'd0;
            10'd229: s <= -16'd10235;
            10'd230: s <= 16'd32433;
            10'd231: s <= -16'd7138;
            10'd232: s <= 16'd4915;
            10'd233: s <= 16'd14936;
            10'd234: s <= -16'd29889;
            10'd235: s <= 16'd6473;
            10'd236: s <= -16'd8514;
            10'd237: s <= -16'd19982;
            10'd238: s <= 16'd25481;
            10'd239: s <= -16'd8421;
            10'd240: s <= 16'd9830;
            10'd241: s <= 16'd24018;
            10'd242: s <= -16'd20394;
            10'd243: s <= 16'd12457;
            10'd244: s <= -16'd8514;
            10'd245: s <= -16'd25966;
            10'd246: s <= 16'd15986;
            10'd247: s <= -16'd17503;
            10'd248: s <= 16'd4915;
            10'd249: s <= 16'd25301;
            10'd250: s <= -16'd13443;
            10'd251: s <= 16'd22203;
            10'd252: s <= 16'd0;
            10'd253: s <= -16'd22204;
            10'd254: s <= 16'd13442;
            10'd255: s <= -16'd25302;
            10'd256: s <= -16'd4916;
            10'd257: s <= 16'd17502;
            10'd258: s <= -16'd15987;
            10'd259: s <= 16'd25965;
            10'd260: s <= 16'd8513;
            10'd261: s <= -16'd12458;
            10'd262: s <= 16'd20393;
            10'd263: s <= -16'd24019;
            10'd264: s <= -16'd9831;
            10'd265: s <= 16'd8420;
            10'd266: s <= -16'd25482;
            10'd267: s <= 16'd19981;
            10'd268: s <= 16'd8513;
            10'd269: s <= -16'd6474;
            10'd270: s <= 16'd29888;
            10'd271: s <= -16'd14937;
            10'd272: s <= -16'd4916;
            10'd273: s <= 16'd7137;
            10'd274: s <= -16'd32434;
            10'd275: s <= 16'd10234;
            10'd276: s <= -16'd1;
            10'd277: s <= -16'd10235;
            10'd278: s <= 16'd32433;
            10'd279: s <= -16'd7138;
            10'd280: s <= 16'd4915;
            10'd281: s <= 16'd14936;
            10'd282: s <= -16'd29889;
            10'd283: s <= 16'd6473;
            10'd284: s <= -16'd8514;
            10'd285: s <= -16'd19982;
            10'd286: s <= 16'd25481;
            10'd287: s <= -16'd8421;
            10'd288: s <= 16'd9830;
            10'd289: s <= 16'd24018;
            10'd290: s <= -16'd20394;
            10'd291: s <= 16'd12457;
            10'd292: s <= -16'd8514;
            10'd293: s <= -16'd25966;
            10'd294: s <= 16'd15986;
            10'd295: s <= -16'd17503;
            10'd296: s <= 16'd4915;
            10'd297: s <= 16'd25301;
            10'd298: s <= -16'd13443;
            10'd299: s <= 16'd22203;
            10'd300: s <= 16'd0;
            10'd301: s <= -16'd22204;
            10'd302: s <= 16'd13442;
            10'd303: s <= -16'd25302;
            10'd304: s <= -16'd4916;
            10'd305: s <= 16'd17502;
            10'd306: s <= -16'd15987;
            10'd307: s <= 16'd25965;
            10'd308: s <= 16'd8513;
            10'd309: s <= -16'd12458;
            10'd310: s <= 16'd20393;
            10'd311: s <= -16'd24019;
            10'd312: s <= -16'd9831;
            10'd313: s <= 16'd8420;
            10'd314: s <= -16'd25482;
            10'd315: s <= 16'd19981;
            10'd316: s <= 16'd8513;
            10'd317: s <= -16'd6474;
            10'd318: s <= 16'd29888;
            10'd319: s <= -16'd14937;
            10'd320: s <= -16'd4916;
            10'd321: s <= 16'd7137;
            10'd322: s <= -16'd32434;
            10'd323: s <= 16'd10234;
            10'd324: s <= -16'd1;
            10'd325: s <= -16'd10235;
            10'd326: s <= 16'd32433;
            10'd327: s <= -16'd7138;
            10'd328: s <= 16'd4915;
            10'd329: s <= 16'd14936;
            10'd330: s <= -16'd29889;
            10'd331: s <= 16'd6473;
            10'd332: s <= -16'd8514;
            10'd333: s <= -16'd19982;
            10'd334: s <= 16'd25481;
            10'd335: s <= -16'd8421;
            10'd336: s <= 16'd9830;
            10'd337: s <= 16'd24018;
            10'd338: s <= -16'd20394;
            10'd339: s <= 16'd12457;
            10'd340: s <= -16'd8514;
            10'd341: s <= -16'd25966;
            10'd342: s <= 16'd15986;
            10'd343: s <= -16'd17503;
            10'd344: s <= 16'd4915;
            10'd345: s <= 16'd25301;
            10'd346: s <= -16'd13443;
            10'd347: s <= 16'd22203;
            10'd348: s <= 16'd0;
            10'd349: s <= -16'd22204;
            10'd350: s <= 16'd13442;
            10'd351: s <= -16'd25302;
            10'd352: s <= -16'd4916;
            10'd353: s <= 16'd17502;
            10'd354: s <= -16'd15987;
            10'd355: s <= 16'd25965;
            10'd356: s <= 16'd8513;
            10'd357: s <= -16'd12458;
            10'd358: s <= 16'd20393;
            10'd359: s <= -16'd24019;
            10'd360: s <= -16'd9831;
            10'd361: s <= 16'd8420;
            10'd362: s <= -16'd25482;
            10'd363: s <= 16'd19981;
            10'd364: s <= 16'd8513;
            10'd365: s <= -16'd6474;
            10'd366: s <= 16'd29888;
            10'd367: s <= -16'd14937;
            10'd368: s <= -16'd4916;
            10'd369: s <= 16'd7137;
            10'd370: s <= -16'd32434;
            10'd371: s <= 16'd10234;
            10'd372: s <= 16'd0;
            10'd373: s <= -16'd10235;
            10'd374: s <= 16'd32433;
            10'd375: s <= -16'd7138;
            10'd376: s <= 16'd4915;
            10'd377: s <= 16'd14936;
            10'd378: s <= -16'd29889;
            10'd379: s <= 16'd6473;
            10'd380: s <= -16'd8514;
            10'd381: s <= -16'd19982;
            10'd382: s <= 16'd25481;
            10'd383: s <= -16'd8421;
            10'd384: s <= 16'd9830;
            10'd385: s <= 16'd24018;
            10'd386: s <= -16'd20394;
            10'd387: s <= 16'd12457;
            10'd388: s <= -16'd8514;
            10'd389: s <= -16'd25966;
            10'd390: s <= 16'd15986;
            10'd391: s <= -16'd17503;
            10'd392: s <= 16'd4915;
            10'd393: s <= 16'd25301;
            10'd394: s <= -16'd13443;
            10'd395: s <= 16'd22203;
            10'd396: s <= -16'd1;
            10'd397: s <= -16'd22204;
            10'd398: s <= 16'd13442;
            10'd399: s <= -16'd25302;
            10'd400: s <= -16'd4916;
            10'd401: s <= 16'd17502;
            10'd402: s <= -16'd15987;
            10'd403: s <= 16'd25965;
            10'd404: s <= 16'd8513;
            10'd405: s <= -16'd12458;
            10'd406: s <= 16'd20393;
            10'd407: s <= -16'd24019;
            10'd408: s <= -16'd9831;
            10'd409: s <= 16'd8420;
            10'd410: s <= -16'd25482;
            10'd411: s <= 16'd19981;
            10'd412: s <= 16'd8513;
            10'd413: s <= -16'd6474;
            10'd414: s <= 16'd29888;
            10'd415: s <= -16'd14937;
            10'd416: s <= -16'd4916;
            10'd417: s <= 16'd7137;
            10'd418: s <= -16'd32434;
            10'd419: s <= 16'd10234;
            10'd420: s <= 16'd0;
            10'd421: s <= -16'd10235;
            10'd422: s <= 16'd32433;
            10'd423: s <= -16'd7138;
            10'd424: s <= 16'd4915;
            10'd425: s <= 16'd14936;
            10'd426: s <= -16'd29889;
            10'd427: s <= 16'd6473;
            10'd428: s <= -16'd8514;
            10'd429: s <= -16'd19982;
            10'd430: s <= 16'd25481;
            10'd431: s <= -16'd8421;
            10'd432: s <= 16'd9830;
            10'd433: s <= 16'd24018;
            10'd434: s <= -16'd20394;
            10'd435: s <= 16'd12457;
            10'd436: s <= -16'd8514;
            10'd437: s <= -16'd25966;
            10'd438: s <= 16'd15986;
            10'd439: s <= -16'd17503;
            10'd440: s <= 16'd4915;
            10'd441: s <= 16'd25301;
            10'd442: s <= -16'd13443;
            10'd443: s <= 16'd22203;
            10'd444: s <= 16'd0;
            10'd445: s <= -16'd22204;
            10'd446: s <= 16'd13442;
            10'd447: s <= -16'd25302;
            10'd448: s <= -16'd4916;
            10'd449: s <= 16'd17502;
            10'd450: s <= -16'd15987;
            10'd451: s <= 16'd25965;
            10'd452: s <= 16'd8513;
            10'd453: s <= -16'd12458;
            10'd454: s <= 16'd20393;
            10'd455: s <= -16'd24019;
            10'd456: s <= -16'd9831;
            10'd457: s <= 16'd8420;
            10'd458: s <= -16'd25482;
            10'd459: s <= 16'd19981;
            10'd460: s <= 16'd8513;
            10'd461: s <= -16'd6474;
            10'd462: s <= 16'd29888;
            10'd463: s <= -16'd14937;
            10'd464: s <= -16'd4916;
            10'd465: s <= 16'd7137;
            10'd466: s <= -16'd32434;
            10'd467: s <= 16'd10234;
            10'd468: s <= 16'd0;
            10'd469: s <= -16'd10235;
            10'd470: s <= 16'd32433;
            10'd471: s <= -16'd7138;
            10'd472: s <= 16'd4915;
            10'd473: s <= 16'd14936;
            10'd474: s <= -16'd29889;
            10'd475: s <= 16'd6473;
            10'd476: s <= -16'd8514;
            10'd477: s <= -16'd19982;
            10'd478: s <= 16'd25481;
            10'd479: s <= -16'd8421;
            10'd480: s <= 16'd9830;
            10'd481: s <= 16'd24018;
            10'd482: s <= -16'd20394;
            10'd483: s <= 16'd12457;
            10'd484: s <= -16'd8514;
            10'd485: s <= -16'd25966;
            10'd486: s <= 16'd15986;
            10'd487: s <= -16'd17503;
            10'd488: s <= 16'd4915;
            10'd489: s <= 16'd25301;
            10'd490: s <= -16'd13443;
            10'd491: s <= 16'd22203;
            10'd492: s <= -16'd1;
            10'd493: s <= -16'd22204;
            10'd494: s <= 16'd13442;
            10'd495: s <= -16'd25302;
            10'd496: s <= -16'd4916;
            10'd497: s <= 16'd17502;
            10'd498: s <= -16'd15987;
            10'd499: s <= 16'd25965;
            10'd500: s <= 16'd8513;
            10'd501: s <= -16'd12458;
            10'd502: s <= 16'd20393;
            10'd503: s <= -16'd24019;
            10'd504: s <= -16'd9831;
            10'd505: s <= 16'd8420;
            10'd506: s <= -16'd25482;
            10'd507: s <= 16'd19981;
            10'd508: s <= 16'd8513;
            10'd509: s <= -16'd6474;
            10'd510: s <= 16'd29888;
            10'd511: s <= -16'd14937;
            10'd512: s <= -16'd4916;
            10'd513: s <= 16'd7137;
            10'd514: s <= -16'd32434;
            10'd515: s <= 16'd10234;
            10'd516: s <= 16'd0;
            10'd517: s <= -16'd10235;
            10'd518: s <= 16'd32433;
            10'd519: s <= -16'd7138;
            10'd520: s <= 16'd4915;
            10'd521: s <= 16'd14936;
            10'd522: s <= -16'd29889;
            10'd523: s <= 16'd6473;
            10'd524: s <= -16'd8514;
            10'd525: s <= -16'd19982;
            10'd526: s <= 16'd25481;
            10'd527: s <= -16'd8421;
            10'd528: s <= 16'd9830;
            10'd529: s <= 16'd24018;
            10'd530: s <= -16'd20394;
            10'd531: s <= 16'd12457;
            10'd532: s <= -16'd8514;
            10'd533: s <= -16'd25966;
            10'd534: s <= 16'd15986;
            10'd535: s <= -16'd17503;
            10'd536: s <= 16'd4915;
            10'd537: s <= 16'd25301;
            10'd538: s <= -16'd13443;
            10'd539: s <= 16'd22203;
            10'd540: s <= -16'd1;
            10'd541: s <= -16'd22204;
            10'd542: s <= 16'd13442;
            10'd543: s <= -16'd25302;
            10'd544: s <= -16'd4916;
            10'd545: s <= 16'd17502;
            10'd546: s <= -16'd15987;
            10'd547: s <= 16'd25965;
            10'd548: s <= 16'd8513;
            10'd549: s <= -16'd12458;
            10'd550: s <= 16'd20393;
            10'd551: s <= -16'd24019;
            10'd552: s <= -16'd9831;
            10'd553: s <= 16'd8420;
            10'd554: s <= -16'd25482;
            10'd555: s <= 16'd19981;
            10'd556: s <= 16'd8513;
            10'd557: s <= -16'd6474;
            10'd558: s <= 16'd29888;
            10'd559: s <= -16'd14937;
            10'd560: s <= -16'd4916;
            10'd561: s <= 16'd7137;
            10'd562: s <= -16'd32434;
            10'd563: s <= 16'd10234;
            10'd564: s <= -16'd1;
            10'd565: s <= -16'd10235;
            10'd566: s <= 16'd32433;
            10'd567: s <= -16'd7138;
            10'd568: s <= 16'd4915;
            10'd569: s <= 16'd14936;
            10'd570: s <= -16'd29889;
            10'd571: s <= 16'd6473;
            10'd572: s <= -16'd8514;
            10'd573: s <= -16'd19982;
            10'd574: s <= 16'd25481;
            10'd575: s <= -16'd8421;
            10'd576: s <= 16'd9830;
            10'd577: s <= 16'd24018;
            10'd578: s <= -16'd20394;
            10'd579: s <= 16'd12457;
            10'd580: s <= -16'd8514;
            10'd581: s <= -16'd25966;
            10'd582: s <= 16'd15986;
            10'd583: s <= -16'd17503;
            10'd584: s <= 16'd4915;
            10'd585: s <= 16'd25301;
            10'd586: s <= -16'd13443;
            10'd587: s <= 16'd22203;
            10'd588: s <= 16'd0;
            10'd589: s <= -16'd22204;
            10'd590: s <= 16'd13442;
            10'd591: s <= -16'd25302;
            10'd592: s <= -16'd4916;
            10'd593: s <= 16'd17502;
            10'd594: s <= -16'd15987;
            10'd595: s <= 16'd25965;
            10'd596: s <= 16'd8513;
            10'd597: s <= -16'd12458;
            10'd598: s <= 16'd20393;
            10'd599: s <= -16'd24019;
            10'd600: s <= -16'd9831;
            10'd601: s <= 16'd8420;
            10'd602: s <= -16'd25482;
            10'd603: s <= 16'd19981;
            10'd604: s <= 16'd8513;
            10'd605: s <= -16'd6474;
            10'd606: s <= 16'd29888;
            10'd607: s <= -16'd14937;
            10'd608: s <= -16'd4916;
            10'd609: s <= 16'd7137;
            10'd610: s <= -16'd32434;
            10'd611: s <= 16'd10234;
            10'd612: s <= 16'd0;
            10'd613: s <= -16'd10235;
            10'd614: s <= 16'd32433;
            10'd615: s <= -16'd7138;
            10'd616: s <= 16'd4915;
            10'd617: s <= 16'd14936;
            10'd618: s <= -16'd29889;
            10'd619: s <= 16'd6473;
            10'd620: s <= -16'd8514;
            10'd621: s <= -16'd19982;
            10'd622: s <= 16'd25481;
            10'd623: s <= -16'd8421;
            10'd624: s <= 16'd9830;
            10'd625: s <= 16'd24018;
            10'd626: s <= -16'd20394;
            10'd627: s <= 16'd12457;
            10'd628: s <= -16'd8514;
            10'd629: s <= -16'd25966;
            10'd630: s <= 16'd15986;
            10'd631: s <= -16'd17503;
            10'd632: s <= 16'd4915;
            10'd633: s <= 16'd25301;
            10'd634: s <= -16'd13443;
            10'd635: s <= 16'd22203;
            10'd636: s <= 16'd0;
            10'd637: s <= -16'd22204;
            10'd638: s <= 16'd13442;
            10'd639: s <= -16'd25302;
            10'd640: s <= -16'd4916;
            10'd641: s <= 16'd17502;
            10'd642: s <= -16'd15987;
            10'd643: s <= 16'd25965;
            10'd644: s <= 16'd8513;
            10'd645: s <= -16'd12458;
            10'd646: s <= 16'd20393;
            10'd647: s <= -16'd24019;
            10'd648: s <= -16'd9831;
            10'd649: s <= 16'd8420;
            10'd650: s <= -16'd25482;
            10'd651: s <= 16'd19981;
            10'd652: s <= 16'd8513;
            10'd653: s <= -16'd6474;
            10'd654: s <= 16'd29888;
            10'd655: s <= -16'd14937;
            10'd656: s <= -16'd4916;
            10'd657: s <= 16'd7137;
            10'd658: s <= -16'd32434;
            10'd659: s <= 16'd10234;
            10'd660: s <= -16'd1;
            10'd661: s <= -16'd10235;
            10'd662: s <= 16'd32433;
            10'd663: s <= -16'd7138;
            10'd664: s <= 16'd4915;
            10'd665: s <= 16'd14936;
            10'd666: s <= -16'd29889;
            10'd667: s <= 16'd6473;
            10'd668: s <= -16'd8514;
            10'd669: s <= -16'd19982;
            10'd670: s <= 16'd25481;
            10'd671: s <= -16'd8421;
            10'd672: s <= 16'd9830;
            10'd673: s <= 16'd24018;
            10'd674: s <= -16'd20394;
            10'd675: s <= 16'd12457;
            10'd676: s <= -16'd8514;
            10'd677: s <= -16'd25966;
            10'd678: s <= 16'd15986;
            10'd679: s <= -16'd17503;
            10'd680: s <= 16'd4915;
            10'd681: s <= 16'd25301;
            10'd682: s <= -16'd13443;
            10'd683: s <= 16'd22203;
            10'd684: s <= 16'd0;
            10'd685: s <= -16'd22204;
            10'd686: s <= 16'd13442;
            10'd687: s <= -16'd25302;
            10'd688: s <= -16'd4916;
            10'd689: s <= 16'd17502;
            10'd690: s <= -16'd15987;
            10'd691: s <= 16'd25965;
            10'd692: s <= 16'd8513;
            10'd693: s <= -16'd12458;
            10'd694: s <= 16'd20393;
            10'd695: s <= -16'd24019;
            10'd696: s <= -16'd9831;
            10'd697: s <= 16'd8420;
            10'd698: s <= -16'd25482;
            10'd699: s <= 16'd19981;
            10'd700: s <= 16'd8513;
            10'd701: s <= -16'd6474;
            10'd702: s <= 16'd29888;
            10'd703: s <= -16'd14937;
            10'd704: s <= -16'd4916;
            10'd705: s <= 16'd7137;
            10'd706: s <= -16'd32434;
            10'd707: s <= 16'd10234;
            10'd708: s <= 16'd0;
            10'd709: s <= -16'd10235;
            10'd710: s <= 16'd32433;
            10'd711: s <= -16'd7138;
            10'd712: s <= 16'd4915;
            10'd713: s <= 16'd14936;
            10'd714: s <= -16'd29889;
            10'd715: s <= 16'd6473;
            10'd716: s <= -16'd8514;
            10'd717: s <= -16'd19982;
            10'd718: s <= 16'd25481;
            10'd719: s <= -16'd8421;
            10'd720: s <= 16'd9830;
            10'd721: s <= 16'd24018;
            10'd722: s <= -16'd20394;
            10'd723: s <= 16'd12457;
            10'd724: s <= -16'd8514;
            10'd725: s <= -16'd25966;
            10'd726: s <= 16'd15986;
            10'd727: s <= -16'd17503;
            10'd728: s <= 16'd4915;
            10'd729: s <= 16'd25301;
            10'd730: s <= -16'd13443;
            10'd731: s <= 16'd22203;
            10'd732: s <= 16'd0;
            10'd733: s <= -16'd22204;
            10'd734: s <= 16'd13442;
            10'd735: s <= -16'd25302;
            10'd736: s <= -16'd4916;
            10'd737: s <= 16'd17502;
            10'd738: s <= -16'd15987;
            10'd739: s <= 16'd25965;
            10'd740: s <= 16'd8513;
            10'd741: s <= -16'd12458;
            10'd742: s <= 16'd20393;
            10'd743: s <= -16'd24019;
            10'd744: s <= -16'd9831;
            10'd745: s <= 16'd8420;
            10'd746: s <= -16'd25482;
            10'd747: s <= 16'd19981;
            10'd748: s <= 16'd8513;
            10'd749: s <= -16'd6474;
            10'd750: s <= 16'd29888;
            10'd751: s <= -16'd14937;
            10'd752: s <= -16'd4916;
            10'd753: s <= 16'd7137;
            10'd754: s <= -16'd32434;
            10'd755: s <= 16'd10234;
            10'd756: s <= -16'd1;
            10'd757: s <= -16'd10235;
            10'd758: s <= 16'd32433;
            10'd759: s <= -16'd7138;
            10'd760: s <= 16'd4915;
            10'd761: s <= 16'd14936;
            10'd762: s <= -16'd29889;
            10'd763: s <= 16'd6473;
            10'd764: s <= -16'd8514;
            10'd765: s <= -16'd19982;
            10'd766: s <= 16'd25481;
            10'd767: s <= -16'd8421;
            10'd768: s <= 16'd9830;
            10'd769: s <= 16'd24018;
            10'd770: s <= -16'd20394;
            10'd771: s <= 16'd12457;
            10'd772: s <= -16'd8514;
            10'd773: s <= -16'd25966;
            10'd774: s <= 16'd15986;
            10'd775: s <= -16'd17503;
            10'd776: s <= 16'd4915;
            10'd777: s <= 16'd25301;
            10'd778: s <= -16'd13443;
            10'd779: s <= 16'd22203;
            10'd780: s <= -16'd1;
            10'd781: s <= -16'd22204;
            10'd782: s <= 16'd13442;
            10'd783: s <= -16'd25302;
            10'd784: s <= -16'd4916;
            10'd785: s <= 16'd17502;
            10'd786: s <= -16'd15987;
            10'd787: s <= 16'd25965;
            10'd788: s <= 16'd8513;
            10'd789: s <= -16'd12458;
            10'd790: s <= 16'd20393;
            10'd791: s <= -16'd24019;
            10'd792: s <= -16'd9831;
            10'd793: s <= 16'd8420;
            10'd794: s <= -16'd25482;
            10'd795: s <= 16'd19981;
            10'd796: s <= 16'd8513;
            10'd797: s <= -16'd6474;
            10'd798: s <= 16'd29888;
            10'd799: s <= -16'd14937;
            10'd800: s <= -16'd4916;
            10'd801: s <= 16'd7137;
            10'd802: s <= -16'd32434;
            10'd803: s <= 16'd10234;
            10'd804: s <= -16'd1;
            10'd805: s <= -16'd10235;
            10'd806: s <= 16'd32433;
            10'd807: s <= -16'd7138;
            10'd808: s <= 16'd4915;
            10'd809: s <= 16'd14936;
            10'd810: s <= -16'd29889;
            10'd811: s <= 16'd6473;
            10'd812: s <= -16'd8514;
            10'd813: s <= -16'd19982;
            10'd814: s <= 16'd25481;
            10'd815: s <= -16'd8421;
            10'd816: s <= 16'd9830;
            10'd817: s <= 16'd24018;
            10'd818: s <= -16'd20394;
            10'd819: s <= 16'd12457;
            10'd820: s <= -16'd8514;
            10'd821: s <= -16'd25966;
            10'd822: s <= 16'd15986;
            10'd823: s <= -16'd17503;
            10'd824: s <= 16'd4915;
            10'd825: s <= 16'd25301;
            10'd826: s <= -16'd13443;
            10'd827: s <= 16'd22203;
            10'd828: s <= 16'd0;
            10'd829: s <= -16'd22204;
            10'd830: s <= 16'd13442;
            10'd831: s <= -16'd25302;
            10'd832: s <= -16'd4916;
            10'd833: s <= 16'd17502;
            10'd834: s <= -16'd15987;
            10'd835: s <= 16'd25965;
            10'd836: s <= 16'd8513;
            10'd837: s <= -16'd12458;
            10'd838: s <= 16'd20393;
            10'd839: s <= -16'd24019;
            10'd840: s <= -16'd9831;
            10'd841: s <= 16'd8420;
            10'd842: s <= -16'd25482;
            10'd843: s <= 16'd19981;
            10'd844: s <= 16'd8513;
            10'd845: s <= -16'd6474;
            10'd846: s <= 16'd29888;
            10'd847: s <= -16'd14937;
            10'd848: s <= -16'd4916;
            10'd849: s <= 16'd7137;
            10'd850: s <= -16'd32434;
            10'd851: s <= 16'd10234;
            10'd852: s <= 16'd0;
            10'd853: s <= -16'd10235;
            10'd854: s <= 16'd32433;
            10'd855: s <= -16'd7138;
            10'd856: s <= 16'd4915;
            10'd857: s <= 16'd14936;
            10'd858: s <= -16'd29889;
            10'd859: s <= 16'd6473;
            10'd860: s <= -16'd8514;
            10'd861: s <= -16'd19982;
            10'd862: s <= 16'd25481;
            10'd863: s <= -16'd8421;
            10'd864: s <= 16'd9830;
            10'd865: s <= 16'd24018;
            10'd866: s <= -16'd20394;
            10'd867: s <= 16'd12457;
            10'd868: s <= -16'd8514;
            10'd869: s <= -16'd25966;
            10'd870: s <= 16'd15986;
            10'd871: s <= -16'd17503;
            10'd872: s <= 16'd4915;
            10'd873: s <= 16'd25301;
            10'd874: s <= -16'd13443;
            10'd875: s <= 16'd22203;
            10'd876: s <= -16'd1;
            10'd877: s <= -16'd22204;
            10'd878: s <= 16'd13442;
            10'd879: s <= -16'd25302;
            10'd880: s <= -16'd4916;
            10'd881: s <= 16'd17502;
            10'd882: s <= -16'd15987;
            10'd883: s <= 16'd25965;
            10'd884: s <= 16'd8513;
            10'd885: s <= -16'd12458;
            10'd886: s <= 16'd20393;
            10'd887: s <= -16'd24019;
            10'd888: s <= -16'd9831;
            10'd889: s <= 16'd8420;
            10'd890: s <= -16'd25482;
            10'd891: s <= 16'd19981;
            10'd892: s <= 16'd8513;
            10'd893: s <= -16'd6474;
            10'd894: s <= 16'd29888;
            10'd895: s <= -16'd14937;
            10'd896: s <= -16'd4916;
            10'd897: s <= 16'd7137;
            10'd898: s <= -16'd32434;
            10'd899: s <= 16'd10234;
            10'd900: s <= -16'd1;
            10'd901: s <= -16'd10235;
            10'd902: s <= 16'd32433;
            10'd903: s <= -16'd7138;
            10'd904: s <= 16'd4915;
            10'd905: s <= 16'd14936;
            10'd906: s <= -16'd29889;
            10'd907: s <= 16'd6473;
            10'd908: s <= -16'd8514;
            10'd909: s <= -16'd19982;
            10'd910: s <= 16'd25481;
            10'd911: s <= -16'd8421;
            10'd912: s <= 16'd9830;
            10'd913: s <= 16'd24018;
            10'd914: s <= -16'd20394;
            10'd915: s <= 16'd12457;
            10'd916: s <= -16'd8514;
            10'd917: s <= -16'd25966;
            10'd918: s <= 16'd15986;
            10'd919: s <= -16'd17503;
            10'd920: s <= 16'd4915;
            10'd921: s <= 16'd25301;
            10'd922: s <= -16'd13443;
            10'd923: s <= 16'd22203;
            10'd924: s <= -16'd1;
            10'd925: s <= -16'd22204;
            10'd926: s <= 16'd13442;
            10'd927: s <= -16'd25302;
            10'd928: s <= -16'd4916;
            10'd929: s <= 16'd17502;
            10'd930: s <= -16'd15987;
            10'd931: s <= 16'd25965;
            10'd932: s <= 16'd8513;
            10'd933: s <= -16'd12458;
            10'd934: s <= 16'd20393;
            10'd935: s <= -16'd24019;
            10'd936: s <= -16'd9831;
            10'd937: s <= 16'd8420;
            10'd938: s <= -16'd25482;
            10'd939: s <= 16'd19981;
            10'd940: s <= 16'd8513;
            10'd941: s <= -16'd6474;
            10'd942: s <= 16'd29888;
            10'd943: s <= -16'd14937;
            10'd944: s <= -16'd4916;
            10'd945: s <= 16'd7137;
            10'd946: s <= -16'd32434;
            10'd947: s <= 16'd10234;
            10'd948: s <= -16'd1;
            10'd949: s <= -16'd10235;
            10'd950: s <= 16'd32433;
            10'd951: s <= -16'd7138;
            10'd952: s <= 16'd4915;
            10'd953: s <= 16'd14936;
            10'd954: s <= -16'd29889;
            10'd955: s <= 16'd6473;
            10'd956: s <= -16'd8514;
            10'd957: s <= -16'd19982;
            10'd958: s <= 16'd25481;
            10'd959: s <= -16'd8421;
            10'd960: s <= 16'd9830;
            10'd961: s <= 16'd24018;
            10'd962: s <= -16'd20394;
            10'd963: s <= 16'd12457;
            10'd964: s <= -16'd8514;
            10'd965: s <= -16'd25966;
            10'd966: s <= 16'd15986;
            10'd967: s <= -16'd17503;
            10'd968: s <= 16'd4915;
            10'd969: s <= 16'd25301;
            10'd970: s <= -16'd13443;
            10'd971: s <= 16'd22203;
            10'd972: s <= -16'd1;
            10'd973: s <= -16'd22204;
            10'd974: s <= 16'd13442;
            10'd975: s <= -16'd25302;
            10'd976: s <= -16'd4916;
            10'd977: s <= 16'd17502;
            10'd978: s <= -16'd15987;
            10'd979: s <= 16'd25965;
            10'd980: s <= 16'd8513;
            10'd981: s <= -16'd12458;
            10'd982: s <= 16'd20393;
            10'd983: s <= -16'd24019;
            10'd984: s <= -16'd9831;
            10'd985: s <= 16'd8420;
            10'd986: s <= -16'd25482;
            10'd987: s <= 16'd19981;
            10'd988: s <= 16'd8513;
            10'd989: s <= -16'd6474;
            10'd990: s <= 16'd29888;
            10'd991: s <= -16'd14937;
            10'd992: s <= -16'd4916;
            10'd993: s <= 16'd7137;
            10'd994: s <= -16'd32434;
            10'd995: s <= 16'd10234;
            10'd996: s <= 16'd0;
            10'd997: s <= -16'd10235;
            10'd998: s <= 16'd32433;
            10'd999: s <= -16'd7138;
            10'd1000: s <= 16'd4915;
            10'd1001: s <= 16'd14936;
            10'd1002: s <= -16'd29889;
            10'd1003: s <= 16'd6473;
            10'd1004: s <= -16'd8514;
            10'd1005: s <= -16'd19982;
            10'd1006: s <= 16'd25481;
            10'd1007: s <= -16'd8421;
            10'd1008: s <= 16'd9830;
            10'd1009: s <= 16'd24018;
            10'd1010: s <= -16'd20394;
            10'd1011: s <= 16'd12457;
            10'd1012: s <= -16'd8514;
            10'd1013: s <= -16'd25966;
            10'd1014: s <= 16'd15986;
            10'd1015: s <= -16'd17503;
            10'd1016: s <= 16'd4915;
            10'd1017: s <= 16'd25301;
            10'd1018: s <= -16'd13443;
            10'd1019: s <= 16'd22203;
            10'd1020: s <= 16'd0;
            10'd1021: s <= -16'd22204;
            10'd1022: s <= 16'd13442;
            10'd1023: s <= -16'd25302;
        endcase
end


endmodule
